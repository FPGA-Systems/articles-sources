--              | |                         |Source code for article 
--==============+=+==============           |"Implementation of the basic components of the DSP Complex multiplier" 
--              | |            ||           |
--    |***|    |***|           ||           |Find more
--====|***|    |***|           \\ |***|     |https://github.com/FPGA-Systems/articles-sources
--====|***|    |***|             =|***|==== |
--====|***|====|***|    |**\                |Read article
--====|***|    |***|====|***\     |***|     |https://fpga-systems.ru/publ/jazyki/vhdl/realizacija_bazovykh_komponentov_cos_kompleksnyj_umnozhitel/4-1-0-131
--    |***|    |***|    |****|====|***|==== |    
--             |***|    |****|    FPGA      |   
--fpga-systems |***| ru |****| developers   |   
--             |***|    |****|  community   |   
--    |***|    |***|    |****|====|***|==== |   
--====|***|    |***|====|***/     |***|     |   
--====|***|====|***|    |**/                |   
--====|***|    |***|             =|***|==== |   
--====|***|    |***|           // |***|     |   
--    |***|    |***|           ||           |   
--              | |            ||           |web      - https://fpga-systems.ru  
--==============+=+==============           |telegram - https://t.me/fpgasystems   
--              | |                         |Youtube  - https://www.youtube.com/c/fpgasystems  

----------------------------------------------------------------------------------------------------------------------------------
-- Author : Vitaly Lotnik
-- Name : complex_multiplier_wrap
-- Created : 23/05/2021
-- v. 0.0.0
----------------------------------------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------------------------------------
-- libraries
----------------------------------------------------------------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library rtl_modem;
    use rtl_modem.pkg_rtl_modem_types.all;

----------------------------------------------------------------------------------------------------------------------------------
-- entity declaration
----------------------------------------------------------------------------------------------------------------------------------
entity complex_multiplier_wrap is
    generic(
          g_a_dw                    : integer := 25
        ; g_b_dw                    : integer := 18
        ; g_type                    : integer := 1
    );
    port(
          iCLK                      : in std_logic
        ; iV                        : in std_logic
        ; iA_I                      : in signed(g_a_dw - 1 downto 0)
        ; iA_Q                      : in signed(g_a_dw - 1 downto 0)
        ; iB_I                      : in signed(g_b_dw - 1 downto 0)
        ; iB_Q                      : in signed(g_b_dw - 1 downto 0)
        ; OV                        : out std_logic
        ; oC_I                      : out signed(g_a_dw + g_b_dw downto 0)
        ; oC_Q                      : out signed(g_a_dw + g_b_dw downto 0)
    );
end;

----------------------------------------------------------------------------------------------------------------------------------
-- architecture declaration
----------------------------------------------------------------------------------------------------------------------------------
architecture behavioral of complex_multiplier_wrap is
----------------------------------------------------------------------------------------------------------------------------------
-- signals declaration
----------------------------------------------------------------------------------------------------------------------------------
    signal ib_v : std_logic;
    signal ib_a : t_iq(i(g_a_dw - 1 downto 0), q(g_a_dw - 1 downto 0));
    signal ib_b : t_iq(i(g_b_dw - 1 downto 0), q(g_b_dw - 1 downto 0));
    signal ob_v : std_logic;
    signal ob_c : t_iq(i(g_a_dw + g_b_dw downto 0), q(g_a_dw + g_b_dw downto 0));

begin
----------------------------------------------------------------------------------------------------------------------------------
-- input
----------------------------------------------------------------------------------------------------------------------------------
    ib_v                            <= iV;
    ib_a.i                          <= iA_I;
    ib_a.q                          <= iA_Q;
    ib_b.i                          <= iB_I;
    ib_b.q                          <= iB_Q;

----------------------------------------------------------------------------------------------------------------------------------
-- connect complex multiplier
----------------------------------------------------------------------------------------------------------------------------------
    u_dsp_cmult : entity rtl_modem.complex_multiplier
    generic map(
          g_a_dw                    => g_a_dw
        , g_b_dw                    => g_b_dw
        , g_type                    => g_type
    )
    port map(
          iCLK                      => iCLK
        , iV                        => ib_v
        , iA                        => ib_a
        , iB                        => ib_b
        , oV                        => ob_v
        , oC                        => ob_c
    );

----------------------------------------------------------------------------------------------------------------------------------
-- output
----------------------------------------------------------------------------------------------------------------------------------
    oV                              <= ob_v;
    oC_I                            <= ob_c.i;
    oC_Q                            <= ob_c.q;

----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------
end;